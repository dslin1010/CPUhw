// Jump_Ctrl

module Jump_Ctrl( Zero,
                  JumpOP
				  // write your code in here
				  );

    input Zero;
	output [1:0] JumpOP;
	// write your code in here
	
endmodule





